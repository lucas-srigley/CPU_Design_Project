module ShiftRight(input wire [31:0] A, B, output wire [31:0] result);
	
	assign result = A >> B;

endmodule