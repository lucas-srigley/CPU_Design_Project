module Encoder_32to5 (output reg [4:0] encoderOutput, input wire [31:0] encoderInput);
    always@(*) 
    begin
		case(encoderInput)
            32'b00000000000000000000000000000001 : encoderOutput <= 5'b00000; //0
            32'b00000000000000000000000000000010 : encoderOutput <= 5'b00001; //1
            32'b00000000000000000000000000000100 : encoderOutput <= 5'b00010; //2
            32'b00000000000000000000000000001000 : encoderOutput <= 5'b00011; //3
            32'b00000000000000000000000000010000 : encoderOutput <= 5'b00100; //4
            32'b00000000000000000000000000100000 : encoderOutput <= 5'b00101; //5
            32'b00000000000000000000000001000000 : encoderOutput <= 5'b00110; //6
            32'b00000000000000000000000010000000 : encoderOutput <= 5'b00111; //7
            32'b00000000000000000000000100000000 : encoderOutput <= 5'b01000; //8
            32'b00000000000000000000001000000000 : encoderOutput <= 5'b01001; //9
            32'b00000000000000000000010000000000 : encoderOutput <= 5'b01010; //10
            32'b00000000000000000000100000000000 : encoderOutput <= 5'b01011; //11
            32'b00000000000000000001000000000000 : encoderOutput <= 5'b01100; //12
            32'b00000000000000000010000000000000 : encoderOutput <= 5'b01101; //13
            32'b00000000000000000100000000000000 : encoderOutput <= 5'b01110; //14
            32'b00000000000000001000000000000000 : encoderOutput <= 5'b01111; //15
            32'b00000000000000010000000000000000 : encoderOutput <= 5'b10000; //16
            32'b00000000000000100000000000000000 : encoderOutput <= 5'b10001; //17
            32'b00000000000001000000000000000000 : encoderOutput <= 5'b10010; //18
            32'b00000000000010000000000000000000 : encoderOutput <= 5'b10011; //19
            32'b00000000000100000000000000000000 : encoderOutput <= 5'b10100; //20
            32'b00000000001000000000000000000000 : encoderOutput <= 5'b10101; //21
            32'b00000000010000000000000000000000 : encoderOutput <= 5'b10110; //22
            32'b00000000100000000000000000000000 : encoderOutput <= 5'b10111; //23
            32'b00000001000000000000000000000000 : encoderOutput <= 5'b11000; //24
            32'b00000010000000000000000000000000 : encoderOutput <= 5'b11001; //25
            32'b00000100000000000000000000000000 : encoderOutput <= 5'b11010; //26
            32'b00001000000000000000000000000000 : encoderOutput <= 5'b11011; //27
            32'b00010000000000000000000000000000 : encoderOutput <= 5'b11100; //28
            32'b00100000000000000000000000000000 : encoderOutput <= 5'b11101; //29
            32'b01000000000000000000000000000000 : encoderOutput <= 5'b11110; //30
            32'b10000000000000000000000000000000 : encoderOutput <= 5'b11111; //31
        endcase
    end
endmodule