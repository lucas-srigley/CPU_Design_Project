module logical_OR (output wire [31:0] result, input wire [31:0] A, B);

	assign result = A | B;

endmodule
