module reg_mdr (
    input wire clear,
    input wire clock,
    input wire enable,
    input wire [31:0] MdataIn,
	 input wire [31:0] BusMuxOut,
    output wire [31:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15
);

endmodule