module SelectEncodeLogic(input [31:0] instr, input wire Gra, Grb, Grc, Rin, Rout, BAout, 
								 output [4:0] opcode, output [31:0] C_sign_extended,
								 output [15:0] RegIn, output [15:0] RegOut);

	 reg [3:0] decoderIn = 4'b0000;
	 reg [15:0] decoderOut;

	 initial
			
	 begin
		RegOut = 16'b0000000000000000;
		RegIn = 16'b0000000000000000;
			 
	 end

	 reg BAout_or_Rout;

	 reg [3:0] RA_GRA, RB_GRB, RC_GRC;

    always@(*)
	 
    begin
	 
    BAout_or_Rout = (Rout | BAout);
	 
    end
	 
	 

    always@(*)
	 
    begin
	 
        RA_GRA = (IR[26:23] & (Gra? 4'b1111: 4'b0000));
        RB_GRB = (IR[22:19] & (Grb? 4'b1111: 4'b0000));
        RC_GRC = (IR[18:15] & (Grc? 4'b1111: 4'b0000));
        decoderIn = (RA_GRA | RB_GRB | RC_GRC );
		  
    end

    always@(*) 
	 
    begin
	 
		case(decoderIn)
            4'b0000 : decoderOut <= 16'b0000000000000001; 
            4'b0001 : decoderOut <= 16'b0000000000000010;
            4'b0010 : decoderOut <= 16'b0000000000000100; 
            4'b0011 : decoderOut <= 16'b0000000000001000; 
            4'b0100 : decoderOut <= 16'b0000000000010000; 
            4'b0101 : decoderOut <= 16'b0000000000100000; 
            4'b0110 : decoderOut <= 16'b0000000001000000;  
            4'b0111 : decoderOut <= 16'b0000000010000000;  
            4'b1000 : decoderOut <= 16'b0000000100000000;  
            4'b1001 : decoderOut <= 16'b0000001000000000;  
            4'b1010 : decoderOut <= 16'b0000010000000000;  
            4'b1011 : decoderOut <= 16'b0000100000000000;  
            4'b1100 : decoderOut <= 16'b0001000000000000;  
            4'b1101 : decoderOut <= 16'b0010000000000000;  
            4'b1110 : decoderOut <= 16'b0100000000000000;  
            4'b1111 : decoderOut <= 16'b1000000000000000; 
			
				// default case
            default: decoderOut  <= 16'b0000000000000000;
				
        endcase
		  
    end

	
	always@(*)
	
    begin
	 
        case(decoderOut)
		  
		  // assign for registers from R0in - R15in
        16'b0000000000000001: RegIn <= 16'b0000000000000001 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000000010: RegIn <= 16'b0000000000000010 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000000100: RegIn <= 16'b0000000000000100 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000001000: RegIn <= 16'b0000000000001000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000010000: RegIn <= 16'b0000000000010000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000100000: RegIn <= 16'b0000000000100000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000001000000: RegIn <= 16'b0000000001000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000010000000: RegIn <= 16'b0000000010000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000100000000: RegIn <= 16'b0000000100000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000001000000000: RegIn <= 16'b0000001000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000010000000000: RegIn <= 16'b0000010000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000100000000000: RegIn <= 16'b0000100000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0001000000000000: RegIn <= 16'b0001000000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0010000000000000: RegIn <= 16'b0010000000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0100000000000000: RegIn <= 16'b0100000000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
        16'b1000000000000000: RegIn <= 16'b1000000000000000 & (Rin ? 16'b1111111111111111: 16'b0000000000000000); 
		  
		  // default case
        default:             RegIn <=  16'b0000000000000000;
		  
        endcase 
		  
    end

   
    always@(*)
	 
    begin
	 
	    case(decoderOut) 
		  
		  // assign for registers from R0out - R15out
        16'b0000000000000001: RegOut <= 16'b0000000000000001 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);
        16'b0000000000000010: RegOut <= 16'b0000000000000010 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);
        16'b0000000000000100: RegOut <= 16'b0000000000000100 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);
        16'b0000000000001000: RegOut <= 16'b0000000000001000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000010000: RegOut <= 16'b0000000000010000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000000100000: RegOut <= 16'b0000000000100000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000); 
        16'b0000000001000000: RegOut <= 16'b0000000001000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0000000010000000: RegOut <= 16'b0000000010000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0000000100000000: RegOut <= 16'b0000000100000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0000001000000000: RegOut <= 16'b0000001000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0000010000000000: RegOut <= 16'b0000010000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0000100000000000: RegOut <= 16'b0000100000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0001000000000000: RegOut <= 16'b0001000000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0010000000000000: RegOut <= 16'b0010000000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b0100000000000000: RegOut <= 16'b0100000000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
        16'b1000000000000000: RegOut <= 16'b1000000000000000 & (BAout_or_Rout? 16'b1111111111111111: 16'b0000000000000000);  
		  
		  // default case
        default:              RegOut <= 16'b0000000000000000;
		  
        endcase 
		  
    end

	always@(instr)
	 
    begin

	    C_sign_extended = $signed(instr[18:0]);

    end
	 
endmodule 
